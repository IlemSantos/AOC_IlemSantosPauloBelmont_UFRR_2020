LIBRARY ieee ;
USE ieee.std_logic_1164.all ;

ENTITY ProcessadorUniciclo IS
	PORT (
	
	);
END ProcessadorUniciclo ;

ARCHITECTURE Behavior OF ProcessadorUniciclo IS

BEGIN

END Behavior ; 